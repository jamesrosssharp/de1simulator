../../hexdriver/hexdriver.vhd